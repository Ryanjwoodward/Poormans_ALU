module palu_bool_logic_unit(input [3:0] a, input [3:0] b, output [3:0] f);

	assign f = a & b;

endmodule